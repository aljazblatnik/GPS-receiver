module TOP (
    input clk,
    input clk2,
    output out,
    output data
);

wire data = clk;

endmodule